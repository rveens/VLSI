`timescale 1ns / 1ps

module fifo_reader #(
    parameter DWIDTH = 32)(
    input clk,
    input rst,
	 output req_in,
    input  ack_in,
    input [0 : DWIDTH-1] data_in,
	 input fifo_empty,
	 output req_out,
    input ack_out,
    output [0 : DWIDTH-1] data_out);
	
    // Output request register
    reg req_out_buf;
    assign req_out = req_out_buf;

    // Input request register
    reg req_in_buf;
    assign req_in = req_in_buf;
	 
    // Accumulator (assigned to output directly)
    reg signed [0:DWIDTH-1] data_out_reg, data_in_reg, temp_data;
    assign data_out = data_in_reg;
	 
	 reg data_ready, temp_flag;
	 
initial begin
    req_in_buf <= 0;
    req_out_buf <= 0;
    data_out_reg <= 0;
	 data_in_reg <= 0;
end
  
    always @(posedge clk) begin
        // Reset => initialize
        if (rst) begin
            req_in_buf <= 0;
            req_out_buf <= 0;
				data_in_reg <= 0;
            data_out_reg <= 0;				
				data_ready <= 0;
        end
        // !Reset => run
        else begin
		  
            // Read handshake complete
            if (req_in && ack_in) begin
					if( !req_out || (req_out && ack_out) ) begin
						data_in_reg <= data_in;	
					end
					else begin
						temp_data <= data_in;
						temp_flag <= 1;
					end
               					
					req_out_buf <= 1;
            end			 

				
			//Read handshake is pending then stop producing output
			if (req_in && !ack_in) begin              
					req_out_buf <= 0;
            end 
								
            // Write handshake complete
            if (req_out && ack_out) begin
					if( temp_flag ) begin
						temp_flag <= 0;
						data_in_reg <= temp_data;
						req_out_buf <= 1;
						req_in_buf <= 1;
					end
              if (fifo_empty == 0) begin
                req_in_buf <= 1;		
              end 
            end 

            //Write handshake is pending then stop acquiring output.
            if (req_out && !ack_out) begin        
					req_in_buf <= 0;
            end 			            			  
				
            // Idle state
            if (!req_in && !ack_in && !req_out && !ack_out) begin
              if (fifo_empty == 0) begin
                req_in_buf <= 1;		
              end			  
            end
				
        end
    end

endmodule
